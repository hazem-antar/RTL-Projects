package cosine_pkg;
  // Function definition as provided earlier
  function signed [7:0] cos_lookup(input signed [7:0] angle);
    case (angle)
      -8'sd128: cos_lookup = 8'sd32;
      -8'sd127: cos_lookup = 8'sd32;
      -8'sd126: cos_lookup = 8'sd32;
      -8'sd125: cos_lookup = 8'sd32;
      -8'sd124: cos_lookup = 8'sd32;
      -8'sd123: cos_lookup = 8'sd32;
      -8'sd122: cos_lookup = 8'sd32;
      -8'sd121: cos_lookup = 8'sd32;
      -8'sd120: cos_lookup = 8'sd31;
      -8'sd119: cos_lookup = 8'sd31;
      -8'sd118: cos_lookup = 8'sd31;
      -8'sd117: cos_lookup = 8'sd31;
      -8'sd116: cos_lookup = 8'sd31;
      -8'sd115: cos_lookup = 8'sd30;
      -8'sd114: cos_lookup = 8'sd30;
      -8'sd113: cos_lookup = 8'sd30;
      -8'sd112: cos_lookup = 8'sd30;
      -8'sd111: cos_lookup = 8'sd29;
      -8'sd110: cos_lookup = 8'sd29;
      -8'sd109: cos_lookup = 8'sd29;
      -8'sd108: cos_lookup = 8'sd28;
      -8'sd107: cos_lookup = 8'sd28;
      -8'sd106: cos_lookup = 8'sd27;
      -8'sd105: cos_lookup = 8'sd27;
      -8'sd104: cos_lookup = 8'sd27;
      -8'sd103: cos_lookup = 8'sd26;
      -8'sd102: cos_lookup = 8'sd26;
      -8'sd101: cos_lookup = 8'sd25;
      -8'sd100: cos_lookup = 8'sd25;
      -8'sd99:  cos_lookup = 8'sd24;
      -8'sd98:  cos_lookup = 8'sd24;
      -8'sd97:  cos_lookup = 8'sd23;
      -8'sd96:  cos_lookup = 8'sd23;
      -8'sd95:  cos_lookup = 8'sd22;
      -8'sd94:  cos_lookup = 8'sd21;
      -8'sd93:  cos_lookup = 8'sd21;
      -8'sd92:  cos_lookup = 8'sd20;
      -8'sd91:  cos_lookup = 8'sd20;
      -8'sd90:  cos_lookup = 8'sd19;
      -8'sd89:  cos_lookup = 8'sd18;
      -8'sd88:  cos_lookup = 8'sd18;
      -8'sd87:  cos_lookup = 8'sd17;
      -8'sd86:  cos_lookup = 8'sd16;
      -8'sd85:  cos_lookup = 8'sd16;
      -8'sd84:  cos_lookup = 8'sd15;
      -8'sd83:  cos_lookup = 8'sd14;
      -8'sd82:  cos_lookup = 8'sd14;
      -8'sd81:  cos_lookup = 8'sd13;
      -8'sd80:  cos_lookup = 8'sd12;
      -8'sd79:  cos_lookup = 8'sd12;
      -8'sd78:  cos_lookup = 8'sd11;
      -8'sd77:  cos_lookup = 8'sd10;
      -8'sd76:  cos_lookup = 8'sd9;
      -8'sd75:  cos_lookup = 8'sd9;
      -8'sd74:  cos_lookup = 8'sd8;
      -8'sd73:  cos_lookup = 8'sd7;
      -8'sd72:  cos_lookup = 8'sd6;
      -8'sd71:  cos_lookup = 8'sd5;
      -8'sd70:  cos_lookup = 8'sd5;
      -8'sd69:  cos_lookup = 8'sd4;
      -8'sd68:  cos_lookup = 8'sd3;
      -8'sd67:  cos_lookup = 8'sd2;
      -8'sd66:  cos_lookup = 8'sd2;
      -8'sd65:  cos_lookup = 8'sd1;
      -8'sd64:  cos_lookup = 8'sd0;
      -8'sd63:  cos_lookup = -8'sd1;
      -8'sd62:  cos_lookup = -8'sd2;
      -8'sd61:  cos_lookup = -8'sd2;
      -8'sd60:  cos_lookup = -8'sd3;
      -8'sd59:  cos_lookup = -8'sd4;
      -8'sd58:  cos_lookup = -8'sd5;
      -8'sd57:  cos_lookup = -8'sd5;
      -8'sd56:  cos_lookup = -8'sd6;
      -8'sd55:  cos_lookup = -8'sd7;
      -8'sd54:  cos_lookup = -8'sd8;
      -8'sd53:  cos_lookup = -8'sd9;
      -8'sd52:  cos_lookup = -8'sd9;
      -8'sd51:  cos_lookup = -8'sd10;
      -8'sd50:  cos_lookup = -8'sd11;
      -8'sd49:  cos_lookup = -8'sd12;
      -8'sd48:  cos_lookup = -8'sd12;
      -8'sd47:  cos_lookup = -8'sd13;
      -8'sd46:  cos_lookup = -8'sd14;
      -8'sd45:  cos_lookup = -8'sd14;
      -8'sd44:  cos_lookup = -8'sd15;
      -8'sd43:  cos_lookup = -8'sd16;
      -8'sd42:  cos_lookup = -8'sd16;
      -8'sd41:  cos_lookup = -8'sd17;
      -8'sd40:  cos_lookup = -8'sd18;
      -8'sd39:  cos_lookup = -8'sd18;
      -8'sd38:  cos_lookup = -8'sd19;
      -8'sd37:  cos_lookup = -8'sd20;
      -8'sd36:  cos_lookup = -8'sd20;
      -8'sd35:  cos_lookup = -8'sd21;
      -8'sd34:  cos_lookup = -8'sd21;
      -8'sd33:  cos_lookup = -8'sd22;
      -8'sd32:  cos_lookup = -8'sd23;
      -8'sd31:  cos_lookup = -8'sd23;
      -8'sd30:  cos_lookup = -8'sd24;
      -8'sd29:  cos_lookup = -8'sd24;
      -8'sd28:  cos_lookup = -8'sd25;
      -8'sd27:  cos_lookup = -8'sd25;
      -8'sd26:  cos_lookup = -8'sd26;
      -8'sd25:  cos_lookup = -8'sd26;
      -8'sd24:  cos_lookup = -8'sd27;
      -8'sd23:  cos_lookup = -8'sd27;
      -8'sd22:  cos_lookup = -8'sd27;
      -8'sd21:  cos_lookup = -8'sd28;
      -8'sd20:  cos_lookup = -8'sd28;
      -8'sd19:  cos_lookup = -8'sd29;
      -8'sd18:  cos_lookup = -8'sd29;
      -8'sd17:  cos_lookup = -8'sd29;
      -8'sd16:  cos_lookup = -8'sd30;
      -8'sd15:  cos_lookup = -8'sd30;
      -8'sd14:  cos_lookup = -8'sd30;
      -8'sd13:  cos_lookup = -8'sd30;
      -8'sd12:  cos_lookup = -8'sd31;
      -8'sd11:  cos_lookup = -8'sd31;
      -8'sd10:  cos_lookup = -8'sd31;
      -8'sd9:   cos_lookup = -8'sd31;
      -8'sd8:   cos_lookup = -8'sd31;
      -8'sd7:   cos_lookup = -8'sd32;
      -8'sd6:   cos_lookup = -8'sd32;
      -8'sd5:   cos_lookup = -8'sd32;
      -8'sd4:   cos_lookup = -8'sd32;
      -8'sd3:   cos_lookup = -8'sd32;
      -8'sd2:   cos_lookup = -8'sd32;
      -8'sd1:   cos_lookup = -8'sd32;
       8'sd0:   cos_lookup = -8'sd32;
       8'sd1:   cos_lookup = -8'sd32;
       8'sd2:   cos_lookup = -8'sd32;
       8'sd3:   cos_lookup = -8'sd32;
       8'sd4:   cos_lookup = -8'sd32;
       8'sd5:   cos_lookup = -8'sd32;
       8'sd6:   cos_lookup = -8'sd32;
       8'sd7:   cos_lookup = -8'sd32;
       8'sd8:   cos_lookup = -8'sd31;
       8'sd9:   cos_lookup = -8'sd31;
       8'sd10:  cos_lookup = -8'sd31;
       8'sd11:  cos_lookup = -8'sd31;
       8'sd12:  cos_lookup = -8'sd31;
       8'sd13:  cos_lookup = -8'sd30;
       8'sd14:  cos_lookup = -8'sd30;
       8'sd15:  cos_lookup = -8'sd30;
       8'sd16:  cos_lookup = -8'sd30;
       8'sd17:  cos_lookup = -8'sd29;
       8'sd18:  cos_lookup = -8'sd29;
       8'sd19:  cos_lookup = -8'sd29;
       8'sd20:  cos_lookup = -8'sd28;
       8'sd21:  cos_lookup = -8'sd28;
       8'sd22:  cos_lookup = -8'sd27;
       8'sd23:  cos_lookup = -8'sd27;
       8'sd24:  cos_lookup = -8'sd27;
       8'sd25:  cos_lookup = -8'sd26;
       8'sd26:  cos_lookup = -8'sd26;
       8'sd27:  cos_lookup = -8'sd25;
       8'sd28:  cos_lookup = -8'sd25;
       8'sd29:  cos_lookup = -8'sd24;
       8'sd30:  cos_lookup = -8'sd24;
       8'sd31:  cos_lookup = -8'sd23;
       8'sd32:  cos_lookup = -8'sd23;
       8'sd33:  cos_lookup = -8'sd22;
       8'sd34:  cos_lookup = -8'sd21;
       8'sd35:  cos_lookup = -8'sd21;
       8'sd36:  cos_lookup = -8'sd20;
       8'sd37:  cos_lookup = -8'sd20;
       8'sd38:  cos_lookup = -8'sd19;
       8'sd39:  cos_lookup = -8'sd18;
       8'sd40:  cos_lookup = -8'sd18;
       8'sd41:  cos_lookup = -8'sd17;
       8'sd42:  cos_lookup = -8'sd16;
       8'sd43:  cos_lookup = -8'sd16;
       8'sd44:  cos_lookup = -8'sd15;
       8'sd45:  cos_lookup = -8'sd14;
       8'sd46:  cos_lookup = -8'sd14;
       8'sd47:  cos_lookup = -8'sd13;
       8'sd48:  cos_lookup = -8'sd12;
       8'sd49:  cos_lookup = -8'sd12;
       8'sd50:  cos_lookup = -8'sd11;
       8'sd51:  cos_lookup = -8'sd10;
       8'sd52:  cos_lookup = -8'sd9;
       8'sd53:  cos_lookup = -8'sd9;
       8'sd54:  cos_lookup = -8'sd8;
       8'sd55:  cos_lookup = -8'sd7;
       8'sd56:  cos_lookup = -8'sd6;
       8'sd57:  cos_lookup = -8'sd5;
       8'sd58:  cos_lookup = -8'sd5;
       8'sd59:  cos_lookup = -8'sd4;
       8'sd60:  cos_lookup = -8'sd3;
       8'sd61:  cos_lookup = -8'sd2;
       8'sd62:  cos_lookup = -8'sd2;
       8'sd63:  cos_lookup = -8'sd1;
       8'sd64:  cos_lookup = 8'sd0;
       8'sd65:  cos_lookup = 8'sd1;
       8'sd66:  cos_lookup = 8'sd2;
       8'sd67:  cos_lookup = 8'sd2;
       8'sd68:  cos_lookup = 8'sd3;
       8'sd69:  cos_lookup = 8'sd4;
       8'sd70:  cos_lookup = 8'sd5;
       8'sd71:  cos_lookup = 8'sd5;
       8'sd72:  cos_lookup = 8'sd6;
       8'sd73:  cos_lookup = 8'sd7;
       8'sd74:  cos_lookup = 8'sd8;
       8'sd75:  cos_lookup = 8'sd9;
       8'sd76:  cos_lookup = 8'sd9;
       8'sd77:  cos_lookup = 8'sd10;
       8'sd78:  cos_lookup = 8'sd11;
       8'sd79:  cos_lookup = 8'sd12;
       8'sd80:  cos_lookup = 8'sd12;
       8'sd81:  cos_lookup = 8'sd13;
       8'sd82:  cos_lookup = 8'sd14;
       8'sd83:  cos_lookup = 8'sd14;
       8'sd84:  cos_lookup = 8'sd15;
       8'sd85:  cos_lookup = 8'sd16;
       8'sd86:  cos_lookup = 8'sd16;
       8'sd87:  cos_lookup = 8'sd17;
       8'sd88:  cos_lookup = 8'sd18;
       8'sd89:  cos_lookup = 8'sd18;
       8'sd90:  cos_lookup = 8'sd19;
       8'sd91:  cos_lookup = 8'sd20;
       8'sd92:  cos_lookup = 8'sd20;
       8'sd93:  cos_lookup = 8'sd21;
       8'sd94:  cos_lookup = 8'sd21;
       8'sd95:  cos_lookup = 8'sd22;
       8'sd96:  cos_lookup = 8'sd23;
       8'sd97:  cos_lookup = 8'sd23;
       8'sd98:  cos_lookup = 8'sd24;
       8'sd99:  cos_lookup = 8'sd24;
       8'sd100: cos_lookup = 8'sd25;
       8'sd101: cos_lookup = 8'sd25;
       8'sd102: cos_lookup = 8'sd26;
       8'sd103: cos_lookup = 8'sd26;
       8'sd104: cos_lookup = 8'sd27;
       8'sd105: cos_lookup = 8'sd27;
       8'sd106: cos_lookup = 8'sd27;
       8'sd107: cos_lookup = 8'sd28;
       8'sd108: cos_lookup = 8'sd28;
       8'sd109: cos_lookup = 8'sd29;
       8'sd110: cos_lookup = 8'sd29;
       8'sd111: cos_lookup = 8'sd29;
       8'sd112: cos_lookup = 8'sd30;
       8'sd113: cos_lookup = 8'sd30;
       8'sd114: cos_lookup = 8'sd30;
       8'sd115: cos_lookup = 8'sd30;
       8'sd116: cos_lookup = 8'sd31;
       8'sd117: cos_lookup = 8'sd31;
       8'sd118: cos_lookup = 8'sd31;
       8'sd119: cos_lookup = 8'sd31;
       8'sd120: cos_lookup = 8'sd31;
       8'sd121: cos_lookup = 8'sd32;
       8'sd122: cos_lookup = 8'sd32;
       8'sd123: cos_lookup = 8'sd32;
       8'sd124: cos_lookup = 8'sd32;
       8'sd125: cos_lookup = 8'sd32;
       8'sd126: cos_lookup = 8'sd32;
       8'sd127: cos_lookup = 8'sd32;
      default:  cos_lookup = 8'sd0; // Default case if necessary
    endcase
	endfunction
endpackage